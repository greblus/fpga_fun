module stupid (input x1, output o);
	assign o = x1;
endmodule