module light (x1, x2, x3, x4, x5, f1, f2, f3, f4, f5, f6, f7, f8);
	input x1, x2, x3, x4, x5;
	output f1, f2, f3, f4, f5, f6, f7, f8;
	assign f1 = x1;
	assign f2 = x2;
	assign f3 = x3;
	assign f4 = x4;
	assign f5 = ~x5;
	assign f6 = ~x5;
	assign f7 = ~x5;
	assign f8 = ~x5;
endmodule